package pkg;
typedef enum logic [2:0] {
  ADD = 3'b000,
  SUB,
  MUL_BIT,
  OR_BIT,
  XOR_BIT,
  NOT,
  LD
} operation;
endpackage


